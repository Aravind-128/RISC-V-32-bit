
`timescale 1ns / 1ps


module pc_adder(
    input [31:0] pc,      // output of program counter is given to this adder
    output [31:0] pc4   );
    
    assign pc4 = pc+4;    // program counter value will be updated
endmodule

